magic
tech sky130A
timestamp 1723631128
<< nwell >>
rect -15 -25 125 190
<< nmos >>
rect 55 -120 70 -70
<< pmos >>
rect 55 -5 70 95
<< ndiff >>
rect 20 -85 55 -70
rect 20 -105 25 -85
rect 45 -105 55 -85
rect 20 -120 55 -105
rect 70 -85 105 -70
rect 70 -105 80 -85
rect 100 -105 105 -85
rect 70 -120 105 -105
<< pdiff >>
rect 20 85 55 95
rect 20 5 25 85
rect 45 5 55 85
rect 20 -5 55 5
rect 70 85 105 95
rect 70 5 80 85
rect 100 5 105 85
rect 70 -5 105 5
<< ndiffc >>
rect 25 -105 45 -85
rect 80 -105 100 -85
<< pdiffc >>
rect 25 5 45 85
rect 80 5 100 85
<< psubdiff >>
rect 5 -160 60 -150
rect 5 -185 20 -160
rect 45 -185 60 -160
rect 5 -195 60 -185
<< nsubdiff >>
rect 5 160 60 170
rect 5 135 20 160
rect 45 135 60 160
rect 5 125 60 135
<< psubdiffcont >>
rect 20 -185 45 -160
<< nsubdiffcont >>
rect 20 135 45 160
<< poly >>
rect 55 95 70 110
rect 55 -25 70 -5
rect 15 -30 70 -25
rect 15 -50 25 -30
rect 45 -50 70 -30
rect 15 -55 70 -50
rect 55 -70 70 -55
rect 55 -135 70 -120
<< polycont >>
rect 25 -50 45 -30
<< locali >>
rect 5 160 60 170
rect 5 135 20 160
rect 45 135 60 160
rect 5 125 60 135
rect 25 95 45 125
rect 20 85 50 95
rect 20 5 25 85
rect 45 5 50 85
rect 20 -5 50 5
rect 75 85 105 95
rect 75 5 80 85
rect 100 5 105 85
rect 75 -5 105 5
rect 80 -25 100 -5
rect 15 -30 55 -25
rect 15 -50 25 -30
rect 45 -50 55 -30
rect 15 -55 55 -50
rect 80 -30 135 -25
rect 80 -50 105 -30
rect 125 -50 135 -30
rect 80 -55 135 -50
rect 25 -85 45 -75
rect 25 -150 45 -105
rect 80 -85 100 -55
rect 80 -115 100 -105
rect 5 -160 60 -150
rect 5 -185 20 -160
rect 45 -185 60 -160
rect 5 -195 60 -185
<< viali >>
rect 20 135 45 160
rect 105 -50 125 -30
rect 20 -185 45 -160
<< metal1 >>
rect 5 160 60 170
rect 5 135 20 160
rect 45 135 60 160
rect 5 125 60 135
rect 80 -30 135 -25
rect 80 -50 105 -30
rect 125 -50 135 -30
rect 80 -55 135 -50
rect 5 -160 60 -150
rect 5 -185 20 -160
rect 45 -185 60 -160
rect 5 -195 60 -185
<< labels >>
rlabel metal1 20 -185 45 -160 1 gnd
rlabel nwell 20 135 45 160 1 Vdd
rlabel viali 105 -50 125 -30 1 Vout
rlabel polycont 25 -50 45 -30 1 Vin
<< end >>
