magic
tech sky130A
timestamp 1724137371
<< nwell >>
rect -60 85 110 180
<< nmos >>
rect 35 0 50 50
<< pmos >>
rect 35 105 50 155
<< ndiff >>
rect 0 35 35 50
rect 0 15 5 35
rect 25 15 35 35
rect 0 0 35 15
rect 50 35 90 50
rect 50 15 60 35
rect 80 15 90 35
rect 50 0 90 15
<< pdiff >>
rect 0 140 35 155
rect 0 120 5 140
rect 25 120 35 140
rect 0 105 35 120
rect 50 140 90 155
rect 50 120 60 140
rect 80 120 90 140
rect 50 105 90 120
<< ndiffc >>
rect 5 15 25 35
rect 60 15 80 35
<< pdiffc >>
rect 5 120 25 140
rect 60 120 80 140
<< psubdiff >>
rect -40 35 0 50
rect -40 15 -35 35
rect -15 15 0 35
rect -40 0 0 15
<< nsubdiff >>
rect -40 140 0 155
rect -40 120 -35 140
rect -15 120 0 140
rect -40 105 0 120
<< psubdiffcont >>
rect -35 15 -15 35
<< nsubdiffcont >>
rect -35 120 -15 140
<< poly >>
rect 35 155 50 170
rect 35 50 50 105
rect 35 -20 50 0
rect -10 -25 50 -20
rect -10 -45 0 -25
rect 25 -45 50 -25
rect -10 -50 50 -45
<< polycont >>
rect 0 -45 25 -25
<< locali >>
rect -40 140 25 150
rect -40 120 -35 140
rect -15 120 5 140
rect -40 105 25 120
rect 5 45 25 105
rect -40 35 25 45
rect -40 15 -35 35
rect -15 15 5 35
rect -40 0 25 15
rect 60 140 80 150
rect 60 35 80 120
rect 60 -20 80 15
rect -60 -25 35 -20
rect -60 -45 0 -25
rect 25 -45 35 -25
rect -60 -50 35 -45
rect 60 -50 110 -20
<< viali >>
rect 5 120 25 140
<< metal1 >>
rect -60 140 110 165
rect -60 120 5 140
rect 25 120 110 140
rect -60 95 110 120
rect -60 -10 110 60
<< labels >>
rlabel locali -60 -30 -60 -30 7 A
port 1 w
rlabel locali 110 -35 110 -35 3 Y
port 2 e
rlabel metal1 -60 130 -60 130 7 Vp
port 3 w
rlabel metal1 -60 20 -60 20 7 Vn
port 4 w
<< end >>
