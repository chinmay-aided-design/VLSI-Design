magic
tech sky130A
timestamp 1724659278
<< nwell >>
rect -65 -20 445 105
<< nmos >>
rect 55 -140 70 -90
rect 255 -140 270 -90
<< pmos >>
rect 55 15 70 65
rect 255 15 270 65
<< ndiff >>
rect 20 -105 55 -90
rect 20 -125 25 -105
rect 45 -125 55 -105
rect 20 -140 55 -125
rect 70 -105 105 -90
rect 70 -125 80 -105
rect 100 -125 105 -105
rect 70 -140 105 -125
rect 220 -105 255 -90
rect 220 -125 225 -105
rect 245 -125 255 -105
rect 220 -140 255 -125
rect 270 -105 305 -90
rect 270 -125 280 -105
rect 300 -125 305 -105
rect 270 -140 305 -125
<< pdiff >>
rect 20 50 55 65
rect 20 30 25 50
rect 45 30 55 50
rect 20 15 55 30
rect 70 50 105 65
rect 70 30 80 50
rect 100 30 105 50
rect 70 15 105 30
rect 220 50 255 65
rect 220 30 225 50
rect 245 30 255 50
rect 220 15 255 30
rect 270 50 305 65
rect 270 30 280 50
rect 300 30 305 50
rect 270 15 305 30
<< ndiffc >>
rect 25 -125 45 -105
rect 80 -125 100 -105
rect 225 -125 245 -105
rect 280 -125 300 -105
<< pdiffc >>
rect 25 30 45 50
rect 80 30 100 50
rect 225 30 245 50
rect 280 30 300 50
<< psubdiff >>
rect 135 -105 190 -95
rect 135 -130 150 -105
rect 175 -130 190 -105
rect 135 -140 190 -130
<< nsubdiff >>
rect -30 50 20 65
rect -30 30 -15 50
rect 5 30 20 50
rect -30 15 20 30
rect 305 50 355 65
rect 305 30 320 50
rect 340 30 355 50
rect 305 15 355 30
<< psubdiffcont >>
rect 150 -130 175 -105
<< nsubdiffcont >>
rect -15 30 5 50
rect 320 30 340 50
<< poly >>
rect 55 65 70 80
rect 255 65 270 80
rect 55 -25 70 15
rect 10 -30 70 -25
rect 10 -50 20 -30
rect 40 -50 70 -30
rect 10 -55 70 -50
rect 55 -90 70 -55
rect 255 -30 270 15
rect 255 -35 315 -30
rect 255 -55 280 -35
rect 300 -55 315 -35
rect 255 -60 315 -55
rect 255 -90 270 -60
rect 55 -155 70 -140
rect 255 -155 270 -140
<< polycont >>
rect 20 -50 40 -30
rect 280 -55 300 -35
<< locali >>
rect -30 50 45 65
rect -30 30 -15 50
rect 5 30 25 50
rect -30 15 45 30
rect 80 50 100 60
rect 80 -25 100 30
rect 220 50 245 65
rect 220 30 225 50
rect 220 -25 245 30
rect 280 50 355 65
rect 300 30 320 50
rect 340 30 355 50
rect 280 15 355 30
rect 10 -30 55 -25
rect 10 -50 20 -30
rect 40 -50 55 -30
rect 10 -55 55 -50
rect 80 -30 245 -25
rect 80 -55 151 -30
rect 176 -55 245 -30
rect 80 -60 245 -55
rect 270 -35 315 -30
rect 270 -55 280 -35
rect 300 -55 315 -35
rect 270 -60 315 -55
rect 25 -105 45 -95
rect 25 -165 45 -125
rect 80 -105 100 -60
rect 80 -135 100 -125
rect 135 -105 190 -95
rect 225 -105 245 -95
rect 135 -130 150 -105
rect 175 -125 225 -105
rect 175 -130 245 -125
rect 135 -140 190 -130
rect 225 -140 245 -130
rect 280 -105 300 -95
rect 280 -165 300 -125
rect 25 -185 300 -165
<< viali >>
rect -15 30 5 50
rect 320 30 340 50
rect 151 -55 176 -30
rect 150 -130 175 -105
<< metal1 >>
rect -30 50 45 65
rect -30 30 -15 50
rect 5 30 45 50
rect -30 15 45 30
rect 220 -25 245 65
rect 280 50 355 65
rect 280 30 320 50
rect 340 30 355 50
rect 280 15 355 30
rect 80 -30 245 -25
rect 80 -55 151 -30
rect 176 -55 245 -30
rect 80 -60 245 -55
rect 135 -105 245 -95
rect 135 -130 150 -105
rect 175 -130 245 -105
rect 135 -140 245 -130
<< labels >>
rlabel locali 20 -30 20 -30 7 A
port 1 w
rlabel locali 280 -35 280 -35 7 B
port 2 w
rlabel metal1 151 -30 151 -30 7 out
port 3 w
rlabel metal1 -15 50 -15 50 7 Vdd
port 4 w
rlabel metal1 340 50 340 50 3 Vdd
port 5 e
rlabel metal1 150 -105 150 -105 7 gnd
port 6 w
<< end >>
