* SPICE3 file created from buf.ext - technology: sky130A


.lib "/usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice" tt

Vpower Vdd gnd 1.8
Vinput Vin gnd PULSE(0 1.8 0 .1n .1n 3n 6.6n 5)


X0 Vout Vin Vdd Vdd sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.35 ps=2.7 w=1 l=0.15
X1 Vout Vin gnd gnd sky130_fd_pr__nfet_01v8 ad=0.175 pd=1.7 as=0.175 ps=1.7 w=0.5 l=0.15

.tran 0.02n 10n
.end
