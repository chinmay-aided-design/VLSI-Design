magic
tech sky130A
timestamp 1724138415
<< locali >>
rect 0 0 20 30
rect 320 0 340 30
<< metal1 >>
rect 0 145 20 215
rect 0 40 20 110
use inv_v3  inv_v3_0
timestamp 1724137371
transform 1 0 60 0 1 50
box -60 -50 110 180
use inv_v3  inv_v3_1
timestamp 1724137371
transform 1 0 230 0 1 50
box -60 -50 110 180
<< labels >>
rlabel metal1 0 180 0 180 7 Vp
rlabel metal1 0 70 0 70 7 Vn
rlabel locali 0 15 0 15 7 Vi
rlabel locali 340 15 340 15 3 Vo
<< end >>
