* SPICE3 file created from buffer.ext - technology: sky130A

X0 inv_v3_1/A Vi Vp Vp sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.175 ps=1.7 w=0.5 l=0.15
X1 inv_v3_1/A Vi Vp Vp sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.175 ps=1.7 w=0.5 l=0.15
X2 Vo inv_v3_1/A Vp Vp sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.75 ps=7 w=0.5 l=0.15
X3 Vo inv_v3_1/A Vp Vp sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.75 ps=7 w=0.5 l=0.15
