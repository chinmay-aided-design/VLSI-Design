magic
tech sky130A
timestamp 1724142645
<< locali >>
rect 0 140 30 170
rect 150 140 170 170
<< metal1 >>
rect 150 140 170 170
rect 290 140 320 170
use inv  inv_0
timestamp 1723631128
transform 1 0 15 0 1 195
box -15 -195 135 190
use inv  inv_1
timestamp 1723631128
transform 1 0 155 0 1 195
box -15 -195 135 190
<< labels >>
rlabel locali 0 155 0 155 7 Vi
port 1 w
rlabel metal1 320 155 320 155 3 Vo
port 2 e
<< end >>
